*Sheet Name:/


* Relay 1
xRelay1 intA +12V intB bit1 GND basicRelay

* Relay 2
xRelay2 intB result intA bit2 GND basicRelay

* Relay 3
xRelay3 overflow intA ignore bit2 GND basicRelay

Vs +12v GND dc 12V ac 0V

*//////////////////////////////////////////////////////////
* Basic Relay using to voltage controlled switches
*//////////////////////////////////////////////////////////
*
* connections:      Normally open terminal
*                   |   Center terminal
*                   |   |   normally closed terminal
*                   |   |   |   positive supply
*                   |   |   |   |   negative supply
*                   |   |   |   |   |
*                   |   |   |   |   |
.subckt basicRelay  1   2   3   4   5

SOpen 1 2 4 5 SW_OPEN on
SClosed 2 3 4 5 SW_CLOSED on

* Some pulldowns, to make sure nothing is floating
R1 1 GND 10k
R2 2 GND 10k
R3 3 GND 10k
R4 4 GND 10k
R5 5 GND 10k

.model SW_OPEN SW(Ron=.1 Roff=1Meg Vt=6 )
.model SW_CLOSED SW(Ron=1Meg Roff=.1 Vt=6 )
.ends

.end
