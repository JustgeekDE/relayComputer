*Sheet Name:/

* Relay 1
xRelay1 +12V OUT GND IN GND basicRelay

* Some pulldowns, to make sure nothing is floating
R1 IN GND 10k
R2 OUT GND 10k

Vs +12v GND dc 12V ac 0V

*//////////////////////////////////////////////////////////
* Basic Relay using to voltage controlled switches
*//////////////////////////////////////////////////////////
*
* connections:      Normally open terminal
*                   |   Center terminal
*                   |   |   normally closed terminal
*                   |   |   |   positive supply
*                   |   |   |   |   negative supply
*                   |   |   |   |   |
*                   |   |   |   |   |
.subckt basicRelay  1   2   3   4   5

SOpen 1 2 4 5 SW_OPEN on
SClosed 2 3 4 5 SW_CLOSED on

.model SW_OPEN SW(Ron=.1 Roff=1Meg Vt=6 )
.model SW_CLOSED SW(Ron=1Meg Roff=.1 Vt=6 )
.ends

.end
